//  @author : Secure, Trusted, and Assured Microelectronics (STAM) Center
//
//  Copyright (c) 2024 STAM Center (SCAI/ASU)
//  Permission is hereby granted, free of charge, to any person obtaining a copy
//  of this software and associated documentation files (the "Software"), to deal
//  in the Software without restriction, including without limitation the rights
//  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
//  copies of the Software, and to permit persons to whom the Software is
//  furnished to do so, subject to the following conditions:
//  The above copyright notice and this permission notice shall be included in
//  all copies or substantial portions of the Software.
//
//  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
//  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
//  THE SOFTWARE.


logic [253:0] test_in_left   = 'h00644e720131a029085045b60181585d07816a910871ca8d0c208c16087cfd46;
logic [253:0] test_in_right  = 'h3058d7e39f03e4a928d7e3a603e4a922d7e3a6f7e4a9228b7e3a6f7ba9228b4a;
logic [253:0] test_key       = 'h265484d5f60a98a1cfd2204308bbcace7939ca61b161a7c3ab5f6495d908c558;
logic [253:0] test_out_left  = 'h284ec006d31aa2caaf108f35c066c62d1d003b50e3686929cf0f8d40929c9dfb;
logic [253:0] test_out_right = 'h1c6ac604dcc0149ee0bb7330cfcc5356a4602559b957b72a822c7a61c75ec6a3;
