//  @author : Secure, Trusted, and Assured Microelectronics (STAM) Center
//
//  Copyright (c) 2024 STAM Center (SCAI/ASU)
//  Permission is hereby granted, free of charge, to any person obtaining a copy
//  of this software and associated documentation files (the "Software"), to deal
//  in the Software without restriction, including without limitation the rights
//  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
//  copies of the Software, and to permit persons to whom the Software is
//  furnished to do so, subject to the following conditions:
//  The above copyright notice and this permission notice shall be included in
//  all copies or substantial portions of the Software.
//
//  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
//  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
//  THE SOFTWARE.


// Module that performs addition between three elements in Galois Field with Prime order
module galois_add_three #(
	parameter N_BITS = 254,
	parameter PRIME_MODULUS = 254'h30644e72e131a029b85045b68181585d2833e84879b9709143e1f593f0000001 // Size: N_BITS
) (
	input  [N_BITS-1:0] num1,
	input  [N_BITS-1:0] num2,
	input  [N_BITS-1:0] num3,
	output [N_BITS-1:0] sum
);

wire [(N_BITS+2)-1:0] temp;
wire signed [(N_BITS+2)-1:0] temp1;
wire signed [(N_BITS+2)-1:0] temp2;

assign temp = num1 + num2 + num3;
assign temp1 = temp - PRIME_MODULUS;
assign temp2 = temp - 2*PRIME_MODULUS;
assign sum = temp2 >= 0 ? temp2[N_BITS-1:0] : temp1 >= 0 ? temp1[N_BITS-1:0] : temp[N_BITS-1:0];

endmodule
